module TLROM( // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185252.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185253.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185254.4]
  output        auto_in_a_ready, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input         auto_in_a_valid, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [2:0]  auto_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [1:0]  auto_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [8:0]  auto_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [16:0] auto_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input  [7:0]  auto_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input         auto_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  input         auto_in_d_ready, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  output        auto_in_d_valid, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  output [1:0]  auto_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  output [8:0]  auto_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
  output [63:0] auto_in_d_bits_data // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185255.4]
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [1:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [8:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [16:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [1:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [8:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
  wire [8:0] index; // @[BootROM.scala 50:34:freechips.rocketchip.system.DefaultFPGAConfig.fir@185816.4]
  wire [3:0] high; // @[BootROM.scala 51:68:freechips.rocketchip.system.DefaultFPGAConfig.fir@185817.4]
  wire  _T_673; // @[BootROM.scala 52:53:freechips.rocketchip.system.DefaultFPGAConfig.fir@185818.4]
  wire [63:0] _GEN_1; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_2; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_3; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_4; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_5; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_6; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_7; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_8; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_9; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_10; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_11; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_12; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_13; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_14; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_15; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_16; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_17; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_18; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_19; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_20; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_21; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_22; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_23; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_24; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_25; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_26; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_27; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_28; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_29; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_30; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_31; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_32; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_33; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_34; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_35; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_36; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_37; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_38; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_39; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_40; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_41; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_42; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_43; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_44; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_45; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_46; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_47; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_48; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_49; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_50; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_51; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_52; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_53; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_54; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_55; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_56; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_57; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_58; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_59; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_60; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_61; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_62; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_63; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_64; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_65; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_66; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_67; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_68; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_69; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_70; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_71; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_72; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_73; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_74; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_75; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_76; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_77; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_78; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_79; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_80; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_81; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_82; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_83; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_84; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_85; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_86; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_87; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_88; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_89; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_90; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_91; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_92; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_93; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_94; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_95; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_96; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_97; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_98; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_99; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_100; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_101; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_102; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_103; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_104; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_105; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_106; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_107; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_108; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_109; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_110; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_111; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_112; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_113; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_114; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_115; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_116; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_117; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_118; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_119; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_120; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_121; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_122; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_123; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_124; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_125; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_126; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_127; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_128; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_129; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_130; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_131; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_132; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_133; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_134; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_135; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_136; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_137; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_138; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_139; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_140; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_141; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_142; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_143; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_144; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_145; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_146; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_147; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_148; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_149; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_150; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_151; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_152; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_153; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_154; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_155; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_156; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_157; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_158; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_159; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_160; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_161; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_162; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_163; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_164; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_165; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_166; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_167; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_168; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_169; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_170; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_171; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_172; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_173; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_174; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_175; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_176; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_177; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_178; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_179; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_180; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_181; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_182; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_183; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_184; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_185; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_186; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_187; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_188; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_189; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_190; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_191; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_192; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_193; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_194; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_195; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_196; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_197; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_198; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_199; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_200; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_201; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_202; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_203; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_204; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_205; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_206; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_207; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_208; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_209; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_210; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_211; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_212; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_213; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_214; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_215; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_216; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_217; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_218; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_219; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_220; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_221; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_222; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_223; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_224; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_225; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_226; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_227; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_228; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_229; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_230; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_231; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_232; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_233; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_234; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_235; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_236; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_237; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_238; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_239; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_240; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_241; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_242; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_243; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_244; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_245; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_246; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_247; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_248; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_249; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_250; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_251; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_252; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_253; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_254; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_255; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_256; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_257; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_258; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_259; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_260; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_261; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_262; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_263; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_264; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_265; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_266; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_267; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_268; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_269; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_270; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_271; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_272; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_273; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_274; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_275; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_276; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_277; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_278; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_279; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_280; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_281; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_282; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_283; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_284; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_285; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_286; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_287; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_288; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_289; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_290; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_291; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_292; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_293; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_294; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_295; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_296; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_297; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_298; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_299; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_300; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_301; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_302; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_303; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_304; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_305; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_306; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_307; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_308; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_309; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_310; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_311; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_312; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_313; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_314; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_315; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_316; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_317; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_318; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_319; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_320; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_321; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_322; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_323; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_324; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_325; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_326; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_327; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_328; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_329; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_330; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_331; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_332; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_333; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_334; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_335; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_336; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_337; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_338; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_339; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_340; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_341; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_342; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_343; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_344; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_345; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_346; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_347; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_348; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_349; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_350; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_351; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_352; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_353; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_354; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_355; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_356; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_357; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_358; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_359; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_360; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_361; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_362; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_363; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_364; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_365; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_366; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_367; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_368; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_369; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_370; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_371; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_372; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_373; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_374; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_375; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_376; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_377; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_378; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_379; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_380; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_381; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_382; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_383; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_384; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_385; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_386; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_387; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_388; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_389; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_390; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_391; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_392; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_393; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_394; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_395; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_396; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_397; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_398; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_399; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_400; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_401; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_402; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_403; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_404; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_405; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_406; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_407; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_408; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_409; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_410; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_411; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_412; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_413; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_414; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_415; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_416; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_417; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_418; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_419; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_420; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_421; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_422; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_423; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_424; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_425; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_426; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_427; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_428; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_429; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_430; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_431; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_432; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_433; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_434; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_435; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_436; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_437; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_438; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_439; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_440; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_441; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_442; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_443; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_444; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_445; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_446; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_447; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_448; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_449; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_450; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_451; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_452; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_453; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_454; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_455; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_456; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_457; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_458; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_459; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_460; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_461; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_462; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_463; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_464; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_465; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_466; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_467; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_468; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_469; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_470; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_471; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_472; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_473; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_474; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_475; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_476; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_477; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_478; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_479; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_480; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_481; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_482; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_483; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_484; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_485; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_486; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_487; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_488; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_489; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_490; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_491; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_492; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_493; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_494; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_495; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_496; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_497; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_498; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_499; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_500; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_501; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_502; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_503; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_504; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_505; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_506; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_507; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_508; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_509; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_510; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  wire [63:0] _GEN_511; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  TLMonitor_41 TLMonitor ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultFPGAConfig.fir@185262.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source)
  );
  assign index = auto_in_a_bits_address[11:3]; // @[BootROM.scala 50:34:freechips.rocketchip.system.DefaultFPGAConfig.fir@185816.4]
  assign high = auto_in_a_bits_address[15:12]; // @[BootROM.scala 51:68:freechips.rocketchip.system.DefaultFPGAConfig.fir@185817.4]
  assign _T_673 = high != 4'h0; // @[BootROM.scala 52:53:freechips.rocketchip.system.DefaultFPGAConfig.fir@185818.4]
  assign _GEN_1 = 9'h1 == index ? 64'h914849b009094b7 : 64'h61000437f1402573; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_2 = 9'h2 == index ? 64'h9094849300c49493 : _GEN_1; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_3 = 9'h3 == index ? 64'h4854849300f49493 : _GEN_2; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_4 = 9'h4 == index ? 64'h8484849300c49493 : _GEN_3; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_5 = 9'h5 == index ? 64'h849b032b34b7e004 : _GEN_4; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_6 = 9'h6 == index ? 64'h849300c49493b2b4 : _GEN_5; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_7 = 9'h7 == index ? 64'h849300c494932b34 : _GEN_6; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_8 = 9'h8 == index ? 64'h849300d49493b2b4 : _GEN_7; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_9 = 9'h9 == index ? 64'hd8e4b7e0045654 : _GEN_8; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_10 = 9'ha == index ? 64'hd494938d94849b : _GEN_9; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_11 = 9'hb == index ? 64'he49493b1b48493 : _GEN_10; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_12 = 9'hc == index ? 64'hc494936c748493 : _GEN_11; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_13 = 9'hd == index ? 64'he4b7e004c6c48493 : _GEN_12; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_14 = 9'he == index ? 64'h94938d94849b00d8 : _GEN_13; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_15 = 9'hf == index ? 64'h9493b1b4849300d4 : _GEN_14; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_16 = 9'h10 == index ? 64'hde070000edfe0dd0 : _GEN_15; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_17 = 9'h11 == index ? 64'h7006000038000000 : _GEN_16; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_18 = 9'h12 == index ? 64'h1100000028000000 : _GEN_17; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_19 = 9'h13 == index ? 64'h10000000 : _GEN_18; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_20 = 9'h14 == index ? 64'h380600006e010000 : _GEN_19; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_21 = 9'h15 == index ? 64'h0 : _GEN_20; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_22 = 9'h16 == index ? 64'h0 : _GEN_21; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_23 = 9'h17 == index ? 64'h1000000 : _GEN_22; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_24 = 9'h18 == index ? 64'h400000003000000 : _GEN_23; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_25 = 9'h19 == index ? 64'h100000000000000 : _GEN_24; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_26 = 9'h1a == index ? 64'h400000003000000 : _GEN_25; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_27 = 9'h1b == index ? 64'h10000000f000000 : _GEN_26; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_28 = 9'h1c == index ? 64'h2100000003000000 : _GEN_27; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_29 = 9'h1d == index ? 64'h656572661b000000 : _GEN_28; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_30 = 9'h1e == index ? 64'h6f722c7370696863 : _GEN_29; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_31 = 9'h1f == index ? 64'h7069686374656b63 : _GEN_30; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_32 = 9'h20 == index ? 64'h6e776f6e6b6e752d : _GEN_31; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_33 = 9'h21 == index ? 64'h7665642d : _GEN_32; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_34 = 9'h22 == index ? 64'h1d00000003000000 : _GEN_33; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_35 = 9'h23 == index ? 64'h6565726626000000 : _GEN_34; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_36 = 9'h24 == index ? 64'h6f722c7370696863 : _GEN_35; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_37 = 9'h25 == index ? 64'h7069686374656b63 : _GEN_36; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_38 = 9'h26 == index ? 64'h6e776f6e6b6e752d : _GEN_37; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_39 = 9'h27 == index ? 64'h100000000000000 : _GEN_38; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_40 = 9'h28 == index ? 64'h73757063 : _GEN_39; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_41 = 9'h29 == index ? 64'h400000003000000 : _GEN_40; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_42 = 9'h2a == index ? 64'h100000000000000 : _GEN_41; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_43 = 9'h2b == index ? 64'h400000003000000 : _GEN_42; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_44 = 9'h2c == index ? 64'hf000000 : _GEN_43; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_45 = 9'h2d == index ? 64'h4075706301000000 : _GEN_44; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_46 = 9'h2e == index ? 64'h300000000000030 : _GEN_45; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_47 = 9'h2f == index ? 64'h2c00000004000000 : _GEN_46; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_48 = 9'h30 == index ? 64'h300000000000000 : _GEN_47; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_49 = 9'h31 == index ? 64'h1b00000015000000 : _GEN_48; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_50 = 9'h32 == index ? 64'h722c657669666973 : _GEN_49; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_51 = 9'h33 == index ? 64'h72003074656b636f : _GEN_50; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_52 = 9'h34 == index ? 64'h76637369 : _GEN_51; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_53 = 9'h35 == index ? 64'h400000003000000 : _GEN_52; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_54 = 9'h36 == index ? 64'h400000003c000000 : _GEN_53; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_55 = 9'h37 == index ? 64'h400000003000000 : _GEN_54; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_56 = 9'h38 == index ? 64'h400000004f000000 : _GEN_55; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_57 = 9'h39 == index ? 64'h400000003000000 : _GEN_56; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_58 = 9'h3a == index ? 64'h1000005c000000 : _GEN_57; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_59 = 9'h3b == index ? 64'h400000003000000 : _GEN_58; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_60 = 9'h3c == index ? 64'h75706369000000 : _GEN_59; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_61 = 9'h3d == index ? 64'h400000003000000 : _GEN_60; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_62 = 9'h3e == index ? 64'h4000000075000000 : _GEN_61; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_63 = 9'h3f == index ? 64'h400000003000000 : _GEN_62; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_64 = 9'h40 == index ? 64'h4000000088000000 : _GEN_63; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_65 = 9'h41 == index ? 64'h400000003000000 : _GEN_64; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_66 = 9'h42 == index ? 64'h10000095000000 : _GEN_65; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_67 = 9'h43 == index ? 64'h400000003000000 : _GEN_66; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_68 = 9'h44 == index ? 64'h1000000a2000000 : _GEN_67; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_69 = 9'h45 == index ? 64'h400000003000000 : _GEN_68; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_70 = 9'h46 == index ? 64'hb3000000 : _GEN_69; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_71 = 9'h47 == index ? 64'h900000003000000 : _GEN_70; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_72 = 9'h48 == index ? 64'h34367672b7000000 : _GEN_71; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_73 = 9'h49 == index ? 64'h63616d69 : _GEN_72; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_74 = 9'h4a == index ? 64'h500000003000000 : _GEN_73; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_75 = 9'h4b == index ? 64'h79616b6fc1000000 : _GEN_74; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_76 = 9'h4c == index ? 64'h300000000000000 : _GEN_75; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_77 = 9'h4d == index ? 64'hc800000004000000 : _GEN_76; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_78 = 9'h4e == index ? 64'h100000040420f00 : _GEN_77; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_79 = 9'h4f == index ? 64'h7075727265746e69 : _GEN_78; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_80 = 9'h50 == index ? 64'h6f72746e6f632d74 : _GEN_79; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_81 = 9'h51 == index ? 64'h72656c6c : _GEN_80; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_82 = 9'h52 == index ? 64'h400000003000000 : _GEN_81; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_83 = 9'h53 == index ? 64'h1000000db000000 : _GEN_82; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_84 = 9'h54 == index ? 64'hf00000003000000 : _GEN_83; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_85 = 9'h55 == index ? 64'h637369721b000000 : _GEN_84; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_86 = 9'h56 == index ? 64'h6e692d7570632c76 : _GEN_85; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_87 = 9'h57 == index ? 64'h300000000006374 : _GEN_86; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_88 = 9'h58 == index ? 64'hec00000000000000 : _GEN_87; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_89 = 9'h59 == index ? 64'h400000003000000 : _GEN_88; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_90 = 9'h5a == index ? 64'h200000001010000 : _GEN_89; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_91 = 9'h5b == index ? 64'h400000003000000 : _GEN_90; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_92 = 9'h5c == index ? 64'h200000007010000 : _GEN_91; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_93 = 9'h5d == index ? 64'h200000002000000 : _GEN_92; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_94 = 9'h5e == index ? 64'h100000002000000 : _GEN_93; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_95 = 9'h5f == index ? 64'h384079726f6d656d : _GEN_94; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_96 = 9'h60 == index ? 64'h30303030303030 : _GEN_95; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_97 = 9'h61 == index ? 64'h700000003000000 : _GEN_96; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_98 = 9'h62 == index ? 64'h6f6d656d69000000 : _GEN_97; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_99 = 9'h63 == index ? 64'h300000000007972 : _GEN_98; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_100 = 9'h64 == index ? 64'hb300000008000000 : _GEN_99; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_101 = 9'h65 == index ? 64'h1000000080 : _GEN_100; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_102 = 9'h66 == index ? 64'h400000003000000 : _GEN_101; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_103 = 9'h67 == index ? 64'h100000001010000 : _GEN_102; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_104 = 9'h68 == index ? 64'h400000003000000 : _GEN_103; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_105 = 9'h69 == index ? 64'h100000007010000 : _GEN_104; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_106 = 9'h6a == index ? 64'h100000002000000 : _GEN_105; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_107 = 9'h6b == index ? 64'h300000000636f73 : _GEN_106; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_108 = 9'h6c == index ? 64'h4000000 : _GEN_107; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_109 = 9'h6d == index ? 64'h300000001000000 : _GEN_108; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_110 = 9'h6e == index ? 64'hf00000004000000 : _GEN_109; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_111 = 9'h6f == index ? 64'h300000001000000 : _GEN_110; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_112 = 9'h70 == index ? 64'h1b0000002c000000 : _GEN_111; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_113 = 9'h71 == index ? 64'h7069686365657266 : _GEN_112; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_114 = 9'h72 == index ? 64'h74656b636f722c73 : _GEN_113; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_115 = 9'h73 == index ? 64'h6b6e752d70696863 : _GEN_114; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_116 = 9'h74 == index ? 64'h636f732d6e776f6e : _GEN_115; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_117 = 9'h75 == index ? 64'h2d656c706d697300 : _GEN_116; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_118 = 9'h76 == index ? 64'h300000000737562 : _GEN_117; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_119 = 9'h77 == index ? 64'hf01000000000000 : _GEN_118; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_120 = 9'h78 == index ? 64'h6e696c6301000000 : _GEN_119; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_121 = 9'h79 == index ? 64'h3030303030324074 : _GEN_120; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_122 = 9'h7a == index ? 64'h300000000000030 : _GEN_121; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_123 = 9'h7b == index ? 64'h1b0000000d000000 : _GEN_122; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_124 = 9'h7c == index ? 64'h6c632c7663736972 : _GEN_123; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_125 = 9'h7d == index ? 64'h30746e69 : _GEN_124; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_126 = 9'h7e == index ? 64'h1000000003000000 : _GEN_125; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_127 = 9'h7f == index ? 64'h200000016010000 : _GEN_126; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_128 = 9'h80 == index ? 64'h200000003000000 : _GEN_127; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_129 = 9'h81 == index ? 64'h300000007000000 : _GEN_128; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_130 = 9'h82 == index ? 64'hb300000008000000 : _GEN_129; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_131 = 9'h83 == index ? 64'h10000000002 : _GEN_130; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_132 = 9'h84 == index ? 64'h800000003000000 : _GEN_131; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_133 = 9'h85 == index ? 64'h746e6f632a010000 : _GEN_132; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_134 = 9'h86 == index ? 64'h2000000006c6f72 : _GEN_133; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_135 = 9'h87 == index ? 64'h7562656401000000 : _GEN_134; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_136 = 9'h88 == index ? 64'h6f72746e6f632d67 : _GEN_135; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_137 = 9'h89 == index ? 64'h304072656c6c : _GEN_136; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_138 = 9'h8a == index ? 64'h2100000003000000 : _GEN_137; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_139 = 9'h8b == index ? 64'h696669731b000000 : _GEN_138; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_140 = 9'h8c == index ? 64'h67756265642c6576 : _GEN_139; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_141 = 9'h8d == index ? 64'h736972003331302d : _GEN_140; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_142 = 9'h8e == index ? 64'h67756265642c7663 : _GEN_141; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_143 = 9'h8f == index ? 64'h3331302d : _GEN_142; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_144 = 9'h90 == index ? 64'h800000003000000 : _GEN_143; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_145 = 9'h91 == index ? 64'h200000016010000 : _GEN_144; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_146 = 9'h92 == index ? 64'h3000000ffff0000 : _GEN_145; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_147 = 9'h93 == index ? 64'hb300000008000000 : _GEN_146; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_148 = 9'h94 == index ? 64'h10000000000000 : _GEN_147; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_149 = 9'h95 == index ? 64'h800000003000000 : _GEN_148; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_150 = 9'h96 == index ? 64'h746e6f632a010000 : _GEN_149; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_151 = 9'h97 == index ? 64'h2000000006c6f72 : _GEN_150; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_152 = 9'h98 == index ? 64'h6f72726501000000 : _GEN_151; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_153 = 9'h99 == index ? 64'h6563697665642d72 : _GEN_152; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_154 = 9'h9a == index ? 64'h3030303340 : _GEN_153; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_155 = 9'h9b == index ? 64'he00000003000000 : _GEN_154; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_156 = 9'h9c == index ? 64'h696669731b000000 : _GEN_155; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_157 = 9'h9d == index ? 64'h726f7272652c6576 : _GEN_156; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_158 = 9'h9e == index ? 64'h300000000000030 : _GEN_157; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_159 = 9'h9f == index ? 64'hb300000008000000 : _GEN_158; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_160 = 9'ha0 == index ? 64'h10000000300000 : _GEN_159; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_161 = 9'ha1 == index ? 64'h100000002000000 : _GEN_160; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_162 = 9'ha2 == index ? 64'h6c616e7265747865 : _GEN_161; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_163 = 9'ha3 == index ? 64'h75727265746e692d : _GEN_162; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_164 = 9'ha4 == index ? 64'h300000000737470 : _GEN_163; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_165 = 9'ha5 == index ? 64'h3401000004000000 : _GEN_164; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_166 = 9'ha6 == index ? 64'h300000003000000 : _GEN_165; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_167 = 9'ha7 == index ? 64'h4501000008000000 : _GEN_166; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_168 = 9'ha8 == index ? 64'h200000001000000 : _GEN_167; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_169 = 9'ha9 == index ? 64'h100000002000000 : _GEN_168; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_170 = 9'haa == index ? 64'h7075727265746e69 : _GEN_169; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_171 = 9'hab == index ? 64'h6f72746e6f632d74 : _GEN_170; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_172 = 9'hac == index ? 64'h3030634072656c6c : _GEN_171; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_173 = 9'had == index ? 64'h30303030 : _GEN_172; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_174 = 9'hae == index ? 64'h400000003000000 : _GEN_173; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_175 = 9'haf == index ? 64'h1000000db000000 : _GEN_174; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_176 = 9'hb0 == index ? 64'hc00000003000000 : _GEN_175; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_177 = 9'hb1 == index ? 64'h637369721b000000 : _GEN_176; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_178 = 9'hb2 == index ? 64'h3063696c702c76 : _GEN_177; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_179 = 9'hb3 == index ? 64'h3000000 : _GEN_178; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_180 = 9'hb4 == index ? 64'h3000000ec000000 : _GEN_179; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_181 = 9'hb5 == index ? 64'h1601000008000000 : _GEN_180; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_182 = 9'hb6 == index ? 64'hb00000002000000 : _GEN_181; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_183 = 9'hb7 == index ? 64'h800000003000000 : _GEN_182; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_184 = 9'hb8 == index ? 64'hcb3000000 : _GEN_183; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_185 = 9'hb9 == index ? 64'h300000000000004 : _GEN_184; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_186 = 9'hba == index ? 64'h2a01000008000000 : _GEN_185; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_187 = 9'hbb == index ? 64'h6c6f72746e6f63 : _GEN_186; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_188 = 9'hbc == index ? 64'h400000003000000 : _GEN_187; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_189 = 9'hbd == index ? 64'h300000050010000 : _GEN_188; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_190 = 9'hbe == index ? 64'h400000003000000 : _GEN_189; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_191 = 9'hbf == index ? 64'h200000063010000 : _GEN_190; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_192 = 9'hc0 == index ? 64'h400000003000000 : _GEN_191; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_193 = 9'hc1 == index ? 64'h300000001010000 : _GEN_192; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_194 = 9'hc2 == index ? 64'h400000003000000 : _GEN_193; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_195 = 9'hc3 == index ? 64'h300000007010000 : _GEN_194; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_196 = 9'hc4 == index ? 64'h100000002000000 : _GEN_195; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_197 = 9'hc5 == index ? 64'h726f702d6f696d6d : _GEN_196; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_198 = 9'hc6 == index ? 64'h3640346978612d74 : _GEN_197; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_199 = 9'hc7 == index ? 64'h30303030303030 : _GEN_198; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_200 = 9'hc8 == index ? 64'h400000003000000 : _GEN_199; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_201 = 9'hc9 == index ? 64'h100000000000000 : _GEN_200; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_202 = 9'hca == index ? 64'h400000003000000 : _GEN_201; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_203 = 9'hcb == index ? 64'h10000000f000000 : _GEN_202; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_204 = 9'hcc == index ? 64'hb00000003000000 : _GEN_203; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_205 = 9'hcd == index ? 64'h706d69731b000000 : _GEN_204; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_206 = 9'hce == index ? 64'h7375622d656c : _GEN_205; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_207 = 9'hcf == index ? 64'hc00000003000000 : _GEN_206; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_208 = 9'hd0 == index ? 64'h600f010000 : _GEN_207; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_209 = 9'hd1 == index ? 64'h2000000060 : _GEN_208; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_210 = 9'hd2 == index ? 64'h100000002000000 : _GEN_209; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_211 = 9'hd3 == index ? 64'h30303031406d6f72 : _GEN_210; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_212 = 9'hd4 == index ? 64'h300000000000030 : _GEN_211; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_213 = 9'hd5 == index ? 64'h1b0000000c000000 : _GEN_212; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_214 = 9'hd6 == index ? 64'h722c657669666973 : _GEN_213; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_215 = 9'hd7 == index ? 64'h300000000306d6f : _GEN_214; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_216 = 9'hd8 == index ? 64'hb300000008000000 : _GEN_215; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_217 = 9'hd9 == index ? 64'h10000000100 : _GEN_216; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_218 = 9'hda == index ? 64'h400000003000000 : _GEN_217; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_219 = 9'hdb == index ? 64'h6d656d2a010000 : _GEN_218; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_220 = 9'hdc == index ? 64'h200000002000000 : _GEN_219; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_221 = 9'hdd == index ? 64'h900000002000000 : _GEN_220; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_222 = 9'hde == index ? 64'h7373657264646123 : _GEN_221; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_223 = 9'hdf == index ? 64'h2300736c6c65632d : _GEN_222; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_224 = 9'he0 == index ? 64'h6c65632d657a6973 : _GEN_223; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_225 = 9'he1 == index ? 64'h61706d6f6300736c : _GEN_224; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_226 = 9'he2 == index ? 64'h6f6d00656c626974 : _GEN_225; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_227 = 9'he3 == index ? 64'h636f6c63006c6564 : _GEN_226; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_228 = 9'he4 == index ? 64'h6575716572662d6b : _GEN_227; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_229 = 9'he5 == index ? 64'h61632d640079636e : _GEN_228; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_230 = 9'he6 == index ? 64'h636f6c622d656863 : _GEN_229; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_231 = 9'he7 == index ? 64'h6400657a69732d6b : _GEN_230; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_232 = 9'he8 == index ? 64'h732d65686361632d : _GEN_231; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_233 = 9'he9 == index ? 64'h61632d6400737465 : _GEN_232; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_234 = 9'hea == index ? 64'h657a69732d656863 : _GEN_233; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_235 = 9'heb == index ? 64'h5f65636976656400 : _GEN_234; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_236 = 9'hec == index ? 64'h632d690065707974 : _GEN_235; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_237 = 9'hed == index ? 64'h6f6c622d65686361 : _GEN_236; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_238 = 9'hee == index ? 64'h657a69732d6b63 : _GEN_237; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_239 = 9'hef == index ? 64'h2d65686361632d69 : _GEN_238; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_240 = 9'hf0 == index ? 64'h632d690073746573 : _GEN_239; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_241 = 9'hf1 == index ? 64'h7a69732d65686361 : _GEN_240; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_242 = 9'hf2 == index ? 64'h6c2d7478656e0065 : _GEN_241; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_243 = 9'hf3 == index ? 64'h6361632d6c657665 : _GEN_242; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_244 = 9'hf4 == index ? 64'h7200676572006568 : _GEN_243; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_245 = 9'hf5 == index ? 64'h6173692c76637369 : _GEN_244; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_246 = 9'hf6 == index ? 64'h73757461747300 : _GEN_245; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_247 = 9'hf7 == index ? 64'h65736162656d6974 : _GEN_246; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_248 = 9'hf8 == index ? 64'h6e6575716572662d : _GEN_247; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_249 = 9'hf9 == index ? 64'h65746e6923007963 : _GEN_248; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_250 = 9'hfa == index ? 64'h65632d7470757272 : _GEN_249; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_251 = 9'hfb == index ? 64'h65746e6900736c6c : _GEN_250; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_252 = 9'hfc == index ? 64'h6f632d7470757272 : _GEN_251; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_253 = 9'hfd == index ? 64'h72656c6c6f72746e : _GEN_252; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_254 = 9'hfe == index ? 64'h702c78756e696c00 : _GEN_253; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_255 = 9'hff == index ? 64'h7200656c646e6168 : _GEN_254; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_256 = 9'h100 == index ? 64'h6e69007365676e61 : _GEN_255; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_257 = 9'h101 == index ? 64'h7374707572726574 : _GEN_256; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_258 = 9'h102 == index ? 64'h65646e657478652d : _GEN_257; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_259 = 9'h103 == index ? 64'h616e2d6765720064 : _GEN_258; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_260 = 9'h104 == index ? 64'h65746e690073656d : _GEN_259; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_261 = 9'h105 == index ? 64'h61702d7470757272 : _GEN_260; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_262 = 9'h106 == index ? 64'h746e6900746e6572 : _GEN_261; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_263 = 9'h107 == index ? 64'h73747075727265 : _GEN_262; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_264 = 9'h108 == index ? 64'h616d2c7663736972 : _GEN_263; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_265 = 9'h109 == index ? 64'h69726f6972702d78 : _GEN_264; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_266 = 9'h10a == index ? 64'h7663736972007974 : _GEN_265; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_267 = 9'h10b == index ? 64'h7665646e2c : _GEN_266; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]  assign _GEN_268 = 9'h10c == index ? 64'h0 : _GEN_267; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_268 = 9'h10c == index ? 64'h0 : _GEN_267; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185835.4]
  assign _GEN_269 = 9'h10d == index ? 64'h0 : _GEN_268; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_270 = 9'h10e == index ? 64'h0 : _GEN_269; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_271 = 9'h10f == index ? 64'h0 : _GEN_270; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_272 = 9'h110 == index ? 64'h0 : _GEN_271; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_273 = 9'h111 == index ? 64'h0 : _GEN_272; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_274 = 9'h112 == index ? 64'h0 : _GEN_273; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_275 = 9'h113 == index ? 64'h0 : _GEN_274; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_276 = 9'h114 == index ? 64'h0 : _GEN_275; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_277 = 9'h115 == index ? 64'h0 : _GEN_276; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_278 = 9'h116 == index ? 64'h0 : _GEN_277; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_279 = 9'h117 == index ? 64'h0 : _GEN_278; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_280 = 9'h118 == index ? 64'h0 : _GEN_279; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_281 = 9'h119 == index ? 64'h0 : _GEN_280; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_282 = 9'h11a == index ? 64'h0 : _GEN_281; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_283 = 9'h11b == index ? 64'h0 : _GEN_282; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_284 = 9'h11c == index ? 64'h0 : _GEN_283; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_285 = 9'h11d == index ? 64'h0 : _GEN_284; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_286 = 9'h11e == index ? 64'h0 : _GEN_285; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_287 = 9'h11f == index ? 64'h0 : _GEN_286; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_288 = 9'h120 == index ? 64'h0 : _GEN_287; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_289 = 9'h121 == index ? 64'h0 : _GEN_288; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_290 = 9'h122 == index ? 64'h0 : _GEN_289; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_291 = 9'h123 == index ? 64'h0 : _GEN_290; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_292 = 9'h124 == index ? 64'h0 : _GEN_291; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_293 = 9'h125 == index ? 64'h0 : _GEN_292; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_294 = 9'h126 == index ? 64'h0 : _GEN_293; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_295 = 9'h127 == index ? 64'h0 : _GEN_294; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_296 = 9'h128 == index ? 64'h0 : _GEN_295; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_297 = 9'h129 == index ? 64'h0 : _GEN_296; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_298 = 9'h12a == index ? 64'h0 : _GEN_297; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_299 = 9'h12b == index ? 64'h0 : _GEN_298; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_300 = 9'h12c == index ? 64'h0 : _GEN_299; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_301 = 9'h12d == index ? 64'h0 : _GEN_300; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_302 = 9'h12e == index ? 64'h0 : _GEN_301; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_303 = 9'h12f == index ? 64'h0 : _GEN_302; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_304 = 9'h130 == index ? 64'h0 : _GEN_303; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_305 = 9'h131 == index ? 64'h0 : _GEN_304; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_306 = 9'h132 == index ? 64'h0 : _GEN_305; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_307 = 9'h133 == index ? 64'h0 : _GEN_306; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_308 = 9'h134 == index ? 64'h0 : _GEN_307; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_309 = 9'h135 == index ? 64'h0 : _GEN_308; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_310 = 9'h136 == index ? 64'h0 : _GEN_309; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_311 = 9'h137 == index ? 64'h0 : _GEN_310; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_312 = 9'h138 == index ? 64'h0 : _GEN_311; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_313 = 9'h139 == index ? 64'h0 : _GEN_312; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_314 = 9'h13a == index ? 64'h0 : _GEN_313; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_315 = 9'h13b == index ? 64'h0 : _GEN_314; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_316 = 9'h13c == index ? 64'h0 : _GEN_315; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_317 = 9'h13d == index ? 64'h0 : _GEN_316; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_318 = 9'h13e == index ? 64'h0 : _GEN_317; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_319 = 9'h13f == index ? 64'h0 : _GEN_318; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_320 = 9'h140 == index ? 64'h0 : _GEN_319; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_321 = 9'h141 == index ? 64'h0 : _GEN_320; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_322 = 9'h142 == index ? 64'h0 : _GEN_321; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_323 = 9'h143 == index ? 64'h0 : _GEN_322; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_324 = 9'h144 == index ? 64'h0 : _GEN_323; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_325 = 9'h145 == index ? 64'h0 : _GEN_324; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_326 = 9'h146 == index ? 64'h0 : _GEN_325; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_327 = 9'h147 == index ? 64'h0 : _GEN_326; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_328 = 9'h148 == index ? 64'h0 : _GEN_327; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_329 = 9'h149 == index ? 64'h0 : _GEN_328; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_330 = 9'h14a == index ? 64'h0 : _GEN_329; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_331 = 9'h14b == index ? 64'h0 : _GEN_330; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_332 = 9'h14c == index ? 64'h0 : _GEN_331; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_333 = 9'h14d == index ? 64'h0 : _GEN_332; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_334 = 9'h14e == index ? 64'h0 : _GEN_333; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_335 = 9'h14f == index ? 64'h0 : _GEN_334; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_336 = 9'h150 == index ? 64'h0 : _GEN_335; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_337 = 9'h151 == index ? 64'h0 : _GEN_336; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_338 = 9'h152 == index ? 64'h0 : _GEN_337; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_339 = 9'h153 == index ? 64'h0 : _GEN_338; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_340 = 9'h154 == index ? 64'h0 : _GEN_339; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_341 = 9'h155 == index ? 64'h0 : _GEN_340; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_342 = 9'h156 == index ? 64'h0 : _GEN_341; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_343 = 9'h157 == index ? 64'h0 : _GEN_342; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_344 = 9'h158 == index ? 64'h0 : _GEN_343; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_345 = 9'h159 == index ? 64'h0 : _GEN_344; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_346 = 9'h15a == index ? 64'h0 : _GEN_345; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_347 = 9'h15b == index ? 64'h0 : _GEN_346; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_348 = 9'h15c == index ? 64'h0 : _GEN_347; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_349 = 9'h15d == index ? 64'h0 : _GEN_348; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_350 = 9'h15e == index ? 64'h0 : _GEN_349; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_351 = 9'h15f == index ? 64'h0 : _GEN_350; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_352 = 9'h160 == index ? 64'h0 : _GEN_351; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_353 = 9'h161 == index ? 64'h0 : _GEN_352; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_354 = 9'h162 == index ? 64'h0 : _GEN_353; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_355 = 9'h163 == index ? 64'h0 : _GEN_354; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_356 = 9'h164 == index ? 64'h0 : _GEN_355; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_357 = 9'h165 == index ? 64'h0 : _GEN_356; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_358 = 9'h166 == index ? 64'h0 : _GEN_357; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_359 = 9'h167 == index ? 64'h0 : _GEN_358; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_360 = 9'h168 == index ? 64'h0 : _GEN_359; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_361 = 9'h169 == index ? 64'h0 : _GEN_360; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_362 = 9'h16a == index ? 64'h0 : _GEN_361; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_363 = 9'h16b == index ? 64'h0 : _GEN_362; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_364 = 9'h16c == index ? 64'h0 : _GEN_363; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_365 = 9'h16d == index ? 64'h0 : _GEN_364; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_366 = 9'h16e == index ? 64'h0 : _GEN_365; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_367 = 9'h16f == index ? 64'h0 : _GEN_366; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_368 = 9'h170 == index ? 64'h0 : _GEN_367; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_369 = 9'h171 == index ? 64'h0 : _GEN_368; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_370 = 9'h172 == index ? 64'h0 : _GEN_369; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_371 = 9'h173 == index ? 64'h0 : _GEN_370; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_372 = 9'h174 == index ? 64'h0 : _GEN_371; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_373 = 9'h175 == index ? 64'h0 : _GEN_372; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_374 = 9'h176 == index ? 64'h0 : _GEN_373; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_375 = 9'h177 == index ? 64'h0 : _GEN_374; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_376 = 9'h178 == index ? 64'h0 : _GEN_375; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_377 = 9'h179 == index ? 64'h0 : _GEN_376; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_378 = 9'h17a == index ? 64'h0 : _GEN_377; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_379 = 9'h17b == index ? 64'h0 : _GEN_378; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_380 = 9'h17c == index ? 64'h0 : _GEN_379; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_381 = 9'h17d == index ? 64'h0 : _GEN_380; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_382 = 9'h17e == index ? 64'h0 : _GEN_381; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_383 = 9'h17f == index ? 64'h0 : _GEN_382; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_384 = 9'h180 == index ? 64'h0 : _GEN_383; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_385 = 9'h181 == index ? 64'h0 : _GEN_384; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_386 = 9'h182 == index ? 64'h0 : _GEN_385; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_387 = 9'h183 == index ? 64'h0 : _GEN_386; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_388 = 9'h184 == index ? 64'h0 : _GEN_387; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_389 = 9'h185 == index ? 64'h0 : _GEN_388; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_390 = 9'h186 == index ? 64'h0 : _GEN_389; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_391 = 9'h187 == index ? 64'h0 : _GEN_390; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_392 = 9'h188 == index ? 64'h0 : _GEN_391; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_393 = 9'h189 == index ? 64'h0 : _GEN_392; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_394 = 9'h18a == index ? 64'h0 : _GEN_393; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_395 = 9'h18b == index ? 64'h0 : _GEN_394; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_396 = 9'h18c == index ? 64'h0 : _GEN_395; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_397 = 9'h18d == index ? 64'h0 : _GEN_396; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_398 = 9'h18e == index ? 64'h0 : _GEN_397; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_399 = 9'h18f == index ? 64'h0 : _GEN_398; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_400 = 9'h190 == index ? 64'h0 : _GEN_399; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_401 = 9'h191 == index ? 64'h0 : _GEN_400; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_402 = 9'h192 == index ? 64'h0 : _GEN_401; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_403 = 9'h193 == index ? 64'h0 : _GEN_402; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_404 = 9'h194 == index ? 64'h0 : _GEN_403; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_405 = 9'h195 == index ? 64'h0 : _GEN_404; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_406 = 9'h196 == index ? 64'h0 : _GEN_405; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_407 = 9'h197 == index ? 64'h0 : _GEN_406; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_408 = 9'h198 == index ? 64'h0 : _GEN_407; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_409 = 9'h199 == index ? 64'h0 : _GEN_408; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_410 = 9'h19a == index ? 64'h0 : _GEN_409; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_411 = 9'h19b == index ? 64'h0 : _GEN_410; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_412 = 9'h19c == index ? 64'h0 : _GEN_411; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_413 = 9'h19d == index ? 64'h0 : _GEN_412; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_414 = 9'h19e == index ? 64'h0 : _GEN_413; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_415 = 9'h19f == index ? 64'h0 : _GEN_414; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_416 = 9'h1a0 == index ? 64'h0 : _GEN_415; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_417 = 9'h1a1 == index ? 64'h0 : _GEN_416; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_418 = 9'h1a2 == index ? 64'h0 : _GEN_417; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_419 = 9'h1a3 == index ? 64'h0 : _GEN_418; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_420 = 9'h1a4 == index ? 64'h0 : _GEN_419; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_421 = 9'h1a5 == index ? 64'h0 : _GEN_420; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_422 = 9'h1a6 == index ? 64'h0 : _GEN_421; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_423 = 9'h1a7 == index ? 64'h0 : _GEN_422; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_424 = 9'h1a8 == index ? 64'h0 : _GEN_423; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_425 = 9'h1a9 == index ? 64'h0 : _GEN_424; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_426 = 9'h1aa == index ? 64'h0 : _GEN_425; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_427 = 9'h1ab == index ? 64'h0 : _GEN_426; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_428 = 9'h1ac == index ? 64'h0 : _GEN_427; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_429 = 9'h1ad == index ? 64'h0 : _GEN_428; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_430 = 9'h1ae == index ? 64'h0 : _GEN_429; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_431 = 9'h1af == index ? 64'h0 : _GEN_430; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_432 = 9'h1b0 == index ? 64'h0 : _GEN_431; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_433 = 9'h1b1 == index ? 64'h0 : _GEN_432; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_434 = 9'h1b2 == index ? 64'h0 : _GEN_433; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_435 = 9'h1b3 == index ? 64'h0 : _GEN_434; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_436 = 9'h1b4 == index ? 64'h0 : _GEN_435; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_437 = 9'h1b5 == index ? 64'h0 : _GEN_436; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_438 = 9'h1b6 == index ? 64'h0 : _GEN_437; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_439 = 9'h1b7 == index ? 64'h0 : _GEN_438; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_440 = 9'h1b8 == index ? 64'h0 : _GEN_439; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_441 = 9'h1b9 == index ? 64'h0 : _GEN_440; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_442 = 9'h1ba == index ? 64'h0 : _GEN_441; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_443 = 9'h1bb == index ? 64'h0 : _GEN_442; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_444 = 9'h1bc == index ? 64'h0 : _GEN_443; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_445 = 9'h1bd == index ? 64'h0 : _GEN_444; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_446 = 9'h1be == index ? 64'h0 : _GEN_445; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_447 = 9'h1bf == index ? 64'h0 : _GEN_446; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_448 = 9'h1c0 == index ? 64'h0 : _GEN_447; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_449 = 9'h1c1 == index ? 64'h0 : _GEN_448; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_450 = 9'h1c2 == index ? 64'h0 : _GEN_449; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_451 = 9'h1c3 == index ? 64'h0 : _GEN_450; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_452 = 9'h1c4 == index ? 64'h0 : _GEN_451; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_453 = 9'h1c5 == index ? 64'h0 : _GEN_452; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_454 = 9'h1c6 == index ? 64'h0 : _GEN_453; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_455 = 9'h1c7 == index ? 64'h0 : _GEN_454; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_456 = 9'h1c8 == index ? 64'h0 : _GEN_455; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_457 = 9'h1c9 == index ? 64'h0 : _GEN_456; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_458 = 9'h1ca == index ? 64'h0 : _GEN_457; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_459 = 9'h1cb == index ? 64'h0 : _GEN_458; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_460 = 9'h1cc == index ? 64'h0 : _GEN_459; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_461 = 9'h1cd == index ? 64'h0 : _GEN_460; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_462 = 9'h1ce == index ? 64'h0 : _GEN_461; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_463 = 9'h1cf == index ? 64'h0 : _GEN_462; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_464 = 9'h1d0 == index ? 64'h0 : _GEN_463; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_465 = 9'h1d1 == index ? 64'h0 : _GEN_464; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_466 = 9'h1d2 == index ? 64'h0 : _GEN_465; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_467 = 9'h1d3 == index ? 64'h0 : _GEN_466; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_468 = 9'h1d4 == index ? 64'h0 : _GEN_467; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_469 = 9'h1d5 == index ? 64'h0 : _GEN_468; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_470 = 9'h1d6 == index ? 64'h0 : _GEN_469; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_471 = 9'h1d7 == index ? 64'h0 : _GEN_470; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_472 = 9'h1d8 == index ? 64'h0 : _GEN_471; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_473 = 9'h1d9 == index ? 64'h0 : _GEN_472; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_474 = 9'h1da == index ? 64'h0 : _GEN_473; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_475 = 9'h1db == index ? 64'h0 : _GEN_474; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_476 = 9'h1dc == index ? 64'h0 : _GEN_475; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_477 = 9'h1dd == index ? 64'h0 : _GEN_476; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_478 = 9'h1de == index ? 64'h0 : _GEN_477; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_479 = 9'h1df == index ? 64'h0 : _GEN_478; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_480 = 9'h1e0 == index ? 64'h0 : _GEN_479; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_481 = 9'h1e1 == index ? 64'h0 : _GEN_480; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_482 = 9'h1e2 == index ? 64'h0 : _GEN_481; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_483 = 9'h1e3 == index ? 64'h0 : _GEN_482; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_484 = 9'h1e4 == index ? 64'h0 : _GEN_483; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_485 = 9'h1e5 == index ? 64'h0 : _GEN_484; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_486 = 9'h1e6 == index ? 64'h0 : _GEN_485; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_487 = 9'h1e7 == index ? 64'h0 : _GEN_486; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_488 = 9'h1e8 == index ? 64'h0 : _GEN_487; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_489 = 9'h1e9 == index ? 64'h0 : _GEN_488; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_490 = 9'h1ea == index ? 64'h0 : _GEN_489; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_491 = 9'h1eb == index ? 64'h0 : _GEN_490; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_492 = 9'h1ec == index ? 64'h0 : _GEN_491; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_493 = 9'h1ed == index ? 64'h0 : _GEN_492; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_494 = 9'h1ee == index ? 64'h0 : _GEN_493; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_495 = 9'h1ef == index ? 64'h0 : _GEN_494; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_496 = 9'h1f0 == index ? 64'h0 : _GEN_495; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_497 = 9'h1f1 == index ? 64'h0 : _GEN_496; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_498 = 9'h1f2 == index ? 64'h0 : _GEN_497; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_499 = 9'h1f3 == index ? 64'h0 : _GEN_498; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_500 = 9'h1f4 == index ? 64'h0 : _GEN_499; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_501 = 9'h1f5 == index ? 64'h0 : _GEN_500; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_502 = 9'h1f6 == index ? 64'h0 : _GEN_501; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_503 = 9'h1f7 == index ? 64'h0 : _GEN_502; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_504 = 9'h1f8 == index ? 64'h0 : _GEN_503; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_505 = 9'h1f9 == index ? 64'h0 : _GEN_504; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_506 = 9'h1fa == index ? 64'h0 : _GEN_505; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_507 = 9'h1fb == index ? 64'h0 : _GEN_506; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_508 = 9'h1fc == index ? 64'h0 : _GEN_507; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_509 = 9'h1fd == index ? 64'h0 : _GEN_508; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_510 = 9'h1fe == index ? 64'h0 : _GEN_509; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign _GEN_511 = 9'h1ff == index ? 64'h0 : _GEN_510; // @[BootROM.scala 52:47:freechips.rocketchip.system.DefaultFPGAConfig.fir@185819.4]
  assign auto_in_a_ready = auto_in_d_ready; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultFPGAConfig.fir@185299.4]
  assign auto_in_d_valid = auto_in_a_valid; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultFPGAConfig.fir@185299.4]
  assign auto_in_d_bits_size = auto_in_a_bits_size; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultFPGAConfig.fir@185299.4]
  assign auto_in_d_bits_source = auto_in_a_bits_source; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultFPGAConfig.fir@185299.4]
  assign auto_in_d_bits_data = _T_673 ? 64'h0 : _GEN_511; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultFPGAConfig.fir@185299.4]
  assign TLMonitor_clock = clock; // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185264.4]
  assign TLMonitor_reset = reset; // @[:freechips.rocketchip.system.DefaultFPGAConfig.fir@185265.4]
  assign TLMonitor_io_in_a_ready = auto_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_d_valid = auto_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_d_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
  assign TLMonitor_io_in_d_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultFPGAConfig.fir@185298.4]
endmodule